module rxtx(clk,
			rst,
			rx,
			tx_vld,
			tx_data,

			rx_vld,
			rx_data,
			tx,
			txrdy);
endmodule
