module regfile(we,
                na,
                nb,
                vn,
                d,
                qa,
                qb);
endmodule
