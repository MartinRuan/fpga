module alu(aluc,
            a,
            b);
endmodule
