module contrl_unit(pc_source,
        aluc,
        wreg,
        );
endmodule
